module descriptor(
input             clk,
input             rst_n,
input             keypoint_valid,
input [31:0]      keypoints,
input             keypoint_done,
input             sobel_valid,
input [15:0]      gradient,
input             channel_x,
input             channel_y,

output            output_valid,
output [31:0]     keypoint,
output [15:0]     descriptor_channel_1,
output [15:0]     descriptor_channel_2,
output [15:0]     descriptor_channel_3,
output [15:0]     descriptor_channel_4,
output            done);

integer count, limit, i, j, k, p, q, r,  o;

reg [31:0] index[0:(N*M)/9];
reg [15:0] grad_intensity[0:((N-2)*(M-2))-1];
reg [15:0] window1[0:15];
reg [15:0] window2[0:15];
reg [15:0] window3[0:15];
reg [15:0] window4[0:15];
reg [15:0] window5[0:15];
reg [15:0] window6[0:15];
reg [15:0] window7[0:15];
reg [15:0] window8[0:15];
reg [15:0] window9[0:15];
reg [15:0] window10[0:15];
reg [15:0] window11[0:15];
reg [15:0] window12[0:15];
reg [15:0] window13[0:15];
reg [15:0] window14[0:15];
reg [15:0] window15[0:15];
reg [15:0] window16[0:15];

reg [15:0] channel1[0:15];
reg [15:0] channel2[0:15];
reg [15:0] channel3[0:15];
reg [15:0] channel4[0:15];

reg [15:0] descriptor_1;
reg [15:0] descriptor_2;
reg [15:0] descriptor_3;
reg [15:0] descriptor_4;

reg [1:0] w1[0:15];
reg [1:0] w2[0:15];
reg [1:0] w3[0:15];
reg [1:0] w4[0:15];
reg [1:0] w5[0:15];
reg [1:0] w6[0:15];
reg [1:0] w7[0:15];
reg [1:0] w8[0:15];
reg [1:0] w9[0:15];
reg [1:0] w10[0:15];
reg [1:0] w11[0:15];
reg [1:0] w12[0:15];
reg [1:0] w13[0:15];
reg [1:0] w14[0:15];
reg [1:0] w15[0:15];
reg [1:0] w16[0:15];

reg [1:0] grad_direction[0:((N-2)*(M-2))-1];
reg [4:0] PS, NS;

parameter IDLE = 4'b0000, GRAD = 4'b0001, ASSIGN = 4'b0010, ROW = 4'b0011, CHECK = 4'b0100, FILL = 4'b0101, PROCESS = 4'b0110, COMPUTE = 4'b0111, KEY = 4'b1000;
parameter N = 450, M = 450;
//parameter N = 480, M = 320;

always @(posedge clk or negedge rst_n)
begin
 if (~rst_n)
  PS <= IDLE;
 else
  PS <= NS;
end

always @(posedge clk)
begin
 if (sobel_valid)
 begin
  grad_intensity[i] <= gradient;
  grad_direction[i] <= (channel_x * 2'b10) + (channel_y * 2'b01);
  i <= (i == ((N-2)*(M-2))-1) ? 0 : i + 1;
 end
 else
  i <= i;
end

always @(posedge clk)
begin
 if (keypoint_valid)
 begin
  index[j] <= keypoints;
  j <= j + 1;
  limit <= j;
 end
 else
 begin
  j <= j;
  limit <= j;
 end
end

always @(sobel_valid, keypoint_valid, keypoint_done, i, count, PS, j, k)
begin
 case (PS)
 IDLE: begin
        i = 0;
        j = 0;
        k = 0;
        o = 0;
        r = 0;
        count = 0;
        if(sobel_valid)
         NS = GRAD;
        else
         NS = IDLE;
       end
 GRAD: begin
        NS = (i == ((N-2)*(M-2))-1) ? KEY : GRAD;
       end
 KEY:  begin
        NS = (keypoint_done == 1) ? ASSIGN : KEY;
       end
 ASSIGN: begin
          o = 0;
          k = index[count];
          count = count + 1;
          NS = (count == limit-1) ? IDLE : ROW;
         end
 ROW: begin
       o = k/M;
       // o = (k-(o*M) > M) ? o + 1 : o;
       NS = (k-(o*M) > M) ? ROW : CHECK;
      end
 CHECK: begin
         NS = (o > 20 && k-(o*M) > 20 && ((o+1)*M)-k > 20 && N-o > 20) ? FILL : ASSIGN;
        end
 FILL: begin
        r = 0;
        for(p = 0; p < 4; p = p+1)
        begin
         for(q = 0; q < 4; q = q+1)
         begin
          window1[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*p)];
          window2[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*p)];
          window3[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*p)];
          window4[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*p)];

          window5[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+4))];
          window6[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+4))];
          window7[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+4))];
          window8[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+4))];

          window9[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+8))];
          window10[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+8))];
          window11[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+8))];
          window12[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+8))];

          window13[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+12))];
          window14[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+12))];
          window15[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+12))];
          window16[r] = grad_intensity[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+12))];

          w1[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*p)];
          w2[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*p)];
          w3[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*p)];
          w4[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*p)];

          w5[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+4))];
          w6[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+4))];
          w7[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+4))];
          w8[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+4))];

          w9[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+8))];
          w10[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+8))];
          w11[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+8))];
          w12[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+8))];

          w13[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + ((M-2)*(p+12))];
          w14[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 4 + ((M-2)*(p+12))];
          w15[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 8 + ((M-2)*(p+12))];
          w16[r] = grad_direction[((k-(M + ((o-1)*2)))-7) + q + 12 + ((M-2)*(p+12))];

          r = r + 1;
         end
        end
        NS = PROCESS;
       end
 PROCESS: begin
           // 00
           channel1[0] = (window1[0]*(~w1[0][1])*(~w1[0][0])) + (window1[1]*(~w1[1][1])*(~w1[1][0])) + (window1[2]*(~w1[2][1])*(~w1[2][0])) + (window1[3]*(~w1[3][1])*(~w1[3][0])) + (window1[4]*(~w1[4][1])*(~w1[4][0])) + (window1[5]*(~w1[5][1])*(~w1[5][0])) + (window1[6]*(~w1[6][1])*(~w1[6][0])) + (window1[7]*(~w1[7][1])*(~w1[7][0])) + (window1[8]*(~w1[8][1])*(~w1[8][0])) + (window1[9]*(~w1[9][1])*(~w1[9][0])) + (window1[10]*(~w1[10][1])*(~w1[10][0])) + (window1[11]*(~w1[11][1])*(~w1[11][0])) +(window1[12]*(~w1[12][1])*(~w1[12][0])) + (window1[13]*(~w1[13][1])*(~w1[13][0])) + (window1[14]*(~w1[14][1])*(~w1[14][0])) + (window1[15]*(~w1[14][1])*(~w1[14][0]));
           // 01
           channel2[0] = (window1[0]*(~w1[0][1])*(w1[0][0])) + (window1[1]*(~w1[1][1])*(w1[1][0])) + (window1[2]*(~w1[2][1])*(w1[2][0])) + (window1[3]*(~w1[3][1])*(w1[3][0])) + (window1[4]*(~w1[4][1])*(w1[4][0])) + (window1[5]*(~w1[5][1])*(w1[5][0])) + (window1[6]*(~w1[6][1])*(w1[6][0])) + (window1[7]*(~w1[7][1])*(w1[7][0])) + (window1[8]*(~w1[8][1])*(w1[8][0])) + (window1[9]*(~w1[9][1])*(w1[9][0])) + (window1[10]*(~w1[10][1])*(w1[10][0])) + (window1[11]*(~w1[11][1])*(w1[11][0])) +(window1[12]*(~w1[12][1])*(w1[12][0])) + (window1[13]*(~w1[13][1])*(w1[13][0])) + (window1[14]*(~w1[14][1])*(w1[14][0])) + (window1[15]*(~w1[14][1])*(w1[14][0]));
           // 10
           channel3[0] = (window1[0]*(w1[0][1])*(~w1[0][0])) + (window1[1]*(w1[1][1])*(~w1[1][0])) + (window1[2]*(w1[2][1])*(~w1[2][0])) + (window1[3]*(w1[3][1])*(~w1[3][0])) + (window1[4]*(w1[4][1])*(~w1[4][0])) + (window1[5]*(w1[5][1])*(~w1[5][0])) + (window1[6]*(w1[6][1])*(~w1[6][0])) + (window1[7]*(w1[7][1])*(~w1[7][0])) + (window1[8]*(w1[8][1])*(~w1[8][0])) + (window1[9]*(w1[9][1])*(~w1[9][0])) + (window1[10]*(w1[10][1])*(~w1[10][0])) + (window1[11]*(w1[11][1])*(~w1[11][0])) +(window1[12]*(w1[12][1])*(~w1[12][0])) + (window1[13]*(w1[13][1])*(~w1[13][0])) + (window1[14]*(w1[14][1])*(~w1[14][0])) + (window1[15]*(w1[14][1])*(~w1[14][0]));
           // 11
           channel4[0] = (window1[0]*(w1[0][1])*(w1[0][0])) + (window1[1]*(w1[1][1])*(w1[1][0])) + (window1[2]*(w1[2][1])*(w1[2][0])) + (window1[3]*(w1[3][1])*(w1[3][0])) + (window1[4]*(w1[4][1])*(w1[4][0])) + (window1[5]*(w1[5][1])*(w1[5][0])) + (window1[6]*(w1[6][1])*(w1[6][0])) + (window1[7]*(w1[7][1])*(w1[7][0])) + (window1[8]*(w1[8][1])*(w1[8][0])) + (window1[9]*(w1[9][1])*(w1[9][0])) + (window1[10]*(w1[10][1])*(w1[10][0])) + (window1[11]*(w1[11][1])*(w1[11][0])) +(window1[12]*(w1[12][1])*(w1[12][0])) + (window1[13]*(w1[13][1])*(w1[13][0])) + (window1[14]*(w1[14][1])*(w1[14][0])) + (window1[15]*(w1[14][1])*(w1[14][0]));

           // 00
           channel1[1] = (window2[0]*(~w2[0][1])*(~w2[0][0])) + (window2[1]*(~w2[1][1])*(~w2[1][0])) + (window2[2]*(~w2[2][1])*(~w2[2][0])) + (window2[3]*(~w2[3][1])*(~w2[3][0])) + (window2[4]*(~w2[4][1])*(~w2[4][0])) + (window2[5]*(~w2[5][1])*(~w2[5][0])) + (window2[6]*(~w2[6][1])*(~w2[6][0])) + (window2[7]*(~w2[7][1])*(~w2[7][0])) + (window2[8]*(~w2[8][1])*(~w2[8][0])) + (window2[9]*(~w2[9][1])*(~w2[9][0])) + (window2[10]*(~w2[10][1])*(~w2[10][0])) + (window2[11]*(~w2[11][1])*(~w2[11][0])) +(window2[12]*(~w2[12][1])*(~w2[12][0])) + (window2[13]*(~w2[13][1])*(~w2[13][0])) + (window2[14]*(~w2[14][1])*(~w2[14][0])) + (window2[15]*(~w2[14][1])*(~w2[14][0]));
           // 01
           channel2[1] = (window2[0]*(~w2[0][1])*(w2[0][0])) + (window2[1]*(~w2[1][1])*(w2[1][0])) + (window2[2]*(~w2[2][1])*(w2[2][0])) + (window2[3]*(~w2[3][1])*(w2[3][0])) + (window2[4]*(~w2[4][1])*(w2[4][0])) + (window2[5]*(~w2[5][1])*(w2[5][0])) + (window2[6]*(~w2[6][1])*(w2[6][0])) + (window2[7]*(~w2[7][1])*(w2[7][0])) + (window2[8]*(~w2[8][1])*(w2[8][0])) + (window2[9]*(~w2[9][1])*(w2[9][0])) + (window2[10]*(~w2[10][1])*(w2[10][0])) + (window2[11]*(~w2[11][1])*(w2[11][0])) +(window2[12]*(~w2[12][1])*(w2[12][0])) + (window2[13]*(~w2[13][1])*(w2[13][0])) + (window2[14]*(~w2[14][1])*(w2[14][0])) + (window2[15]*(~w2[14][1])*(w2[14][0]));
           // 10
           channel3[1] = (window2[0]*(w2[0][1])*(~w2[0][0])) + (window2[1]*(w2[1][1])*(~w2[1][0])) + (window2[2]*(w2[2][1])*(~w2[2][0])) + (window2[3]*(w2[3][1])*(~w2[3][0])) + (window2[4]*(w2[4][1])*(~w2[4][0])) + (window2[5]*(w2[5][1])*(~w2[5][0])) + (window2[6]*(w2[6][1])*(~w2[6][0])) + (window2[7]*(w2[7][1])*(~w2[7][0])) + (window2[8]*(w2[8][1])*(~w2[8][0])) + (window2[9]*(w2[9][1])*(~w2[9][0])) + (window2[10]*(w2[10][1])*(~w2[10][0])) + (window2[11]*(w2[11][1])*(~w2[11][0])) +(window2[12]*(w2[12][1])*(~w2[12][0])) + (window2[13]*(w2[13][1])*(~w2[13][0])) + (window2[14]*(w2[14][1])*(~w2[14][0])) + (window2[15]*(w2[14][1])*(~w2[14][0]));
           // 11
           channel4[1] = (window2[0]*(w2[0][1])*(w2[0][0])) + (window2[1]*(w2[1][1])*(w2[1][0])) + (window2[2]*(w2[2][1])*(w2[2][0])) + (window2[3]*(w2[3][1])*(w2[3][0])) + (window2[4]*(w2[4][1])*(w2[4][0])) + (window2[5]*(w2[5][1])*(w2[5][0])) + (window2[6]*(w2[6][1])*(w2[6][0])) + (window2[7]*(w2[7][1])*(w2[7][0])) + (window2[8]*(w2[8][1])*(w2[8][0])) + (window2[9]*(w2[9][1])*(w2[9][0])) + (window2[10]*(w2[10][1])*(w2[10][0])) + (window2[11]*(w2[11][1])*(w2[11][0])) +(window2[12]*(w2[12][1])*(w2[12][0])) + (window2[13]*(w2[13][1])*(w2[13][0])) + (window2[14]*(w2[14][1])*(w2[14][0])) + (window2[15]*(w2[14][1])*(w2[14][0]));

           // 00
           channel1[2] = (window3[0]*(~w3[0][1])*(~w3[0][0])) + (window3[1]*(~w3[1][1])*(~w3[1][0])) + (window3[2]*(~w3[2][1])*(~w3[2][0])) + (window3[3]*(~w3[3][1])*(~w3[3][0])) + (window3[4]*(~w3[4][1])*(~w3[4][0])) + (window3[5]*(~w3[5][1])*(~w3[5][0])) + (window3[6]*(~w3[6][1])*(~w3[6][0])) + (window3[7]*(~w3[7][1])*(~w3[7][0])) + (window3[8]*(~w3[8][1])*(~w3[8][0])) + (window3[9]*(~w3[9][1])*(~w3[9][0])) + (window3[10]*(~w3[10][1])*(~w3[10][0])) + (window3[11]*(~w3[11][1])*(~w3[11][0])) +(window3[12]*(~w3[12][1])*(~w3[12][0])) + (window3[13]*(~w3[13][1])*(~w3[13][0])) + (window3[14]*(~w3[14][1])*(~w3[14][0])) + (window3[15]*(~w3[14][1])*(~w3[14][0]));
           // 01
           channel2[2] = (window3[0]*(~w3[0][1])*(w3[0][0])) + (window3[1]*(~w3[1][1])*(w3[1][0])) + (window3[2]*(~w3[2][1])*(w3[2][0])) + (window3[3]*(~w3[3][1])*(w3[3][0])) + (window3[4]*(~w3[4][1])*(w3[4][0])) + (window3[5]*(~w3[5][1])*(w3[5][0])) + (window3[6]*(~w3[6][1])*(w3[6][0])) + (window3[7]*(~w3[7][1])*(w3[7][0])) + (window3[8]*(~w3[8][1])*(w3[8][0])) + (window3[9]*(~w3[9][1])*(w3[9][0])) + (window3[10]*(~w3[10][1])*(w3[10][0])) + (window3[11]*(~w3[11][1])*(w3[11][0])) +(window3[12]*(~w3[12][1])*(w3[12][0])) + (window3[13]*(~w3[13][1])*(w3[13][0])) + (window3[14]*(~w3[14][1])*(w3[14][0])) + (window3[15]*(~w3[14][1])*(w3[14][0]));
           // 10
           channel3[2] = (window3[0]*(w3[0][1])*(~w3[0][0])) + (window3[1]*(w3[1][1])*(~w3[1][0])) + (window3[2]*(w3[2][1])*(~w3[2][0])) + (window3[3]*(w3[3][1])*(~w3[3][0])) + (window3[4]*(w3[4][1])*(~w3[4][0])) + (window3[5]*(w3[5][1])*(~w3[5][0])) + (window3[6]*(w3[6][1])*(~w3[6][0])) + (window3[7]*(w3[7][1])*(~w3[7][0])) + (window3[8]*(w3[8][1])*(~w3[8][0])) + (window3[9]*(w3[9][1])*(~w3[9][0])) + (window3[10]*(w3[10][1])*(~w3[10][0])) + (window3[11]*(w3[11][1])*(~w3[11][0])) +(window3[12]*(w3[12][1])*(~w3[12][0])) + (window3[13]*(w3[13][1])*(~w3[13][0])) + (window3[14]*(w3[14][1])*(~w3[14][0])) + (window3[15]*(w3[14][1])*(~w3[14][0]));
           // 11
           channel4[2] = (window3[0]*(w3[0][1])*(w3[0][0])) + (window3[1]*(w3[1][1])*(w3[1][0])) + (window3[2]*(w3[2][1])*(w3[2][0])) + (window3[3]*(w3[3][1])*(w3[3][0])) + (window3[4]*(w3[4][1])*(w3[4][0])) + (window3[5]*(w3[5][1])*(w3[5][0])) + (window3[6]*(w3[6][1])*(w3[6][0])) + (window3[7]*(w3[7][1])*(w3[7][0])) + (window3[8]*(w3[8][1])*(w3[8][0])) + (window3[9]*(w3[9][1])*(w3[9][0])) + (window3[10]*(w3[10][1])*(w3[10][0])) + (window3[11]*(w3[11][1])*(w3[11][0])) +(window3[12]*(w3[12][1])*(w3[12][0])) + (window3[13]*(w3[13][1])*(w3[13][0])) + (window3[14]*(w3[14][1])*(w3[14][0])) + (window3[15]*(w3[14][1])*(w3[14][0]));

           // 00
           channel1[3] = (window4[0]*(~w4[0][1])*(~w4[0][0])) + (window4[1]*(~w4[1][1])*(~w4[1][0])) + (window4[2]*(~w4[2][1])*(~w4[2][0])) + (window4[3]*(~w4[3][1])*(~w4[3][0])) + (window4[4]*(~w4[4][1])*(~w4[4][0])) + (window4[5]*(~w4[5][1])*(~w4[5][0])) + (window4[6]*(~w4[6][1])*(~w4[6][0])) + (window4[7]*(~w4[7][1])*(~w4[7][0])) + (window4[8]*(~w4[8][1])*(~w4[8][0])) + (window4[9]*(~w4[9][1])*(~w4[9][0])) + (window4[10]*(~w4[10][1])*(~w4[10][0])) + (window4[11]*(~w4[11][1])*(~w4[11][0])) +(window4[12]*(~w4[12][1])*(~w4[12][0])) + (window4[13]*(~w4[13][1])*(~w4[13][0])) + (window4[14]*(~w4[14][1])*(~w4[14][0])) + (window4[15]*(~w4[14][1])*(~w4[14][0]));
           // 01
           channel2[3] = (window4[0]*(~w4[0][1])*(w4[0][0])) + (window4[1]*(~w4[1][1])*(w4[1][0])) + (window4[2]*(~w4[2][1])*(w4[2][0])) + (window4[3]*(~w4[3][1])*(w4[3][0])) + (window4[4]*(~w4[4][1])*(w4[4][0])) + (window4[5]*(~w4[5][1])*(w4[5][0])) + (window4[6]*(~w4[6][1])*(w4[6][0])) + (window4[7]*(~w4[7][1])*(w4[7][0])) + (window4[8]*(~w4[8][1])*(w4[8][0])) + (window4[9]*(~w4[9][1])*(w4[9][0])) + (window4[10]*(~w4[10][1])*(w4[10][0])) + (window4[11]*(~w4[11][1])*(w4[11][0])) +(window4[12]*(~w4[12][1])*(w4[12][0])) + (window4[13]*(~w4[13][1])*(w4[13][0])) + (window4[14]*(~w4[14][1])*(w4[14][0])) + (window4[15]*(~w4[14][1])*(w4[14][0]));
           // 10
           channel3[3] = (window4[0]*(w4[0][1])*(~w4[0][0])) + (window4[1]*(w4[1][1])*(~w4[1][0])) + (window4[2]*(w4[2][1])*(~w4[2][0])) + (window4[3]*(w4[3][1])*(~w4[3][0])) + (window4[4]*(w4[4][1])*(~w4[4][0])) + (window4[5]*(w4[5][1])*(~w4[5][0])) + (window4[6]*(w4[6][1])*(~w4[6][0])) + (window4[7]*(w4[7][1])*(~w4[7][0])) + (window4[8]*(w4[8][1])*(~w4[8][0])) + (window4[9]*(w4[9][1])*(~w4[9][0])) + (window4[10]*(w4[10][1])*(~w4[10][0])) + (window4[11]*(w4[11][1])*(~w4[11][0])) +(window4[12]*(w4[12][1])*(~w4[12][0])) + (window4[13]*(w4[13][1])*(~w4[13][0])) + (window4[14]*(w4[14][1])*(~w4[14][0])) + (window4[15]*(w4[14][1])*(~w4[14][0]));
           // 11
           channel4[3] = (window4[0]*(w4[0][1])*(w4[0][0])) + (window4[1]*(w4[1][1])*(w4[1][0])) + (window4[2]*(w4[2][1])*(w4[2][0])) + (window4[3]*(w4[3][1])*(w4[3][0])) + (window4[4]*(w4[4][1])*(w4[4][0])) + (window4[5]*(w4[5][1])*(w4[5][0])) + (window4[6]*(w4[6][1])*(w4[6][0])) + (window4[7]*(w4[7][1])*(w4[7][0])) + (window4[8]*(w4[8][1])*(w4[8][0])) + (window4[9]*(w4[9][1])*(w4[9][0])) + (window4[10]*(w4[10][1])*(w4[10][0])) + (window4[11]*(w4[11][1])*(w4[11][0])) +(window4[12]*(w4[12][1])*(w4[12][0])) + (window4[13]*(w4[13][1])*(w4[13][0])) + (window4[14]*(w4[14][1])*(w4[14][0])) + (window4[15]*(w4[14][1])*(w4[14][0]));

           // 00
           channel1[4] = (window5[0]*(~w5[0][1])*(~w5[0][0])) + (window5[1]*(~w5[1][1])*(~w5[1][0])) + (window5[2]*(~w5[2][1])*(~w5[2][0])) + (window5[3]*(~w5[3][1])*(~w5[3][0])) + (window5[4]*(~w5[4][1])*(~w5[4][0])) + (window5[5]*(~w5[5][1])*(~w5[5][0])) + (window5[6]*(~w5[6][1])*(~w5[6][0])) + (window5[7]*(~w5[7][1])*(~w5[7][0])) + (window5[8]*(~w5[8][1])*(~w5[8][0])) + (window5[9]*(~w5[9][1])*(~w5[9][0])) + (window5[10]*(~w5[10][1])*(~w5[10][0])) + (window5[11]*(~w5[11][1])*(~w5[11][0])) +(window5[12]*(~w5[12][1])*(~w5[12][0])) + (window5[13]*(~w5[13][1])*(~w5[13][0])) + (window5[14]*(~w5[14][1])*(~w5[14][0])) + (window5[15]*(~w5[14][1])*(~w5[14][0]));
           // 01
           channel2[4] = (window5[0]*(~w5[0][1])*(w5[0][0])) + (window5[1]*(~w5[1][1])*(w5[1][0])) + (window5[2]*(~w5[2][1])*(w5[2][0])) + (window5[3]*(~w5[3][1])*(w5[3][0])) + (window5[4]*(~w5[4][1])*(w5[4][0])) + (window5[5]*(~w5[5][1])*(w5[5][0])) + (window5[6]*(~w5[6][1])*(w5[6][0])) + (window5[7]*(~w5[7][1])*(w5[7][0])) + (window5[8]*(~w5[8][1])*(w5[8][0])) + (window5[9]*(~w5[9][1])*(w5[9][0])) + (window5[10]*(~w5[10][1])*(w5[10][0])) + (window5[11]*(~w5[11][1])*(w5[11][0])) +(window5[12]*(~w5[12][1])*(w5[12][0])) + (window5[13]*(~w5[13][1])*(w5[13][0])) + (window5[14]*(~w5[14][1])*(w5[14][0])) + (window5[15]*(~w5[14][1])*(w5[14][0]));
           // 10
           channel3[4] = (window5[0]*(w5[0][1])*(~w5[0][0])) + (window5[1]*(w5[1][1])*(~w5[1][0])) + (window5[2]*(w5[2][1])*(~w5[2][0])) + (window5[3]*(w5[3][1])*(~w5[3][0])) + (window5[4]*(w5[4][1])*(~w5[4][0])) + (window5[5]*(w5[5][1])*(~w5[5][0])) + (window5[6]*(w5[6][1])*(~w5[6][0])) + (window5[7]*(w5[7][1])*(~w5[7][0])) + (window5[8]*(w5[8][1])*(~w5[8][0])) + (window5[9]*(w5[9][1])*(~w5[9][0])) + (window5[10]*(w5[10][1])*(~w5[10][0])) + (window5[11]*(w5[11][1])*(~w5[11][0])) +(window5[12]*(w5[12][1])*(~w5[12][0])) + (window5[13]*(w5[13][1])*(~w5[13][0])) + (window5[14]*(w5[14][1])*(~w5[14][0])) + (window5[15]*(w5[14][1])*(~w5[14][0]));
           // 11
           channel4[4] = (window5[0]*(w5[0][1])*(w5[0][0])) + (window5[1]*(w5[1][1])*(w5[1][0])) + (window5[2]*(w5[2][1])*(w5[2][0])) + (window5[3]*(w5[3][1])*(w5[3][0])) + (window5[4]*(w5[4][1])*(w5[4][0])) + (window5[5]*(w5[5][1])*(w5[5][0])) + (window5[6]*(w5[6][1])*(w5[6][0])) + (window5[7]*(w5[7][1])*(w5[7][0])) + (window5[8]*(w5[8][1])*(w5[8][0])) + (window5[9]*(w5[9][1])*(w5[9][0])) + (window5[10]*(w5[10][1])*(w5[10][0])) + (window5[11]*(w5[11][1])*(w5[11][0])) +(window5[12]*(w5[12][1])*(w5[12][0])) + (window5[13]*(w5[13][1])*(w5[13][0])) + (window5[14]*(w5[14][1])*(w5[14][0])) + (window5[15]*(w5[14][1])*(w5[14][0]));

           // 00
           channel1[5] = (window6[0]*(~w6[0][1])*(~w6[0][0])) + (window6[1]*(~w6[1][1])*(~w6[1][0])) + (window6[2]*(~w6[2][1])*(~w6[2][0])) + (window6[3]*(~w6[3][1])*(~w6[3][0])) + (window6[4]*(~w6[4][1])*(~w6[4][0])) + (window6[5]*(~w6[5][1])*(~w6[5][0])) + (window6[6]*(~w6[6][1])*(~w6[6][0])) + (window6[7]*(~w6[7][1])*(~w6[7][0])) + (window6[8]*(~w6[8][1])*(~w6[8][0])) + (window6[9]*(~w6[9][1])*(~w6[9][0])) + (window6[10]*(~w6[10][1])*(~w6[10][0])) + (window6[11]*(~w6[11][1])*(~w6[11][0])) +(window6[12]*(~w6[12][1])*(~w6[12][0])) + (window6[13]*(~w6[13][1])*(~w6[13][0])) + (window6[14]*(~w6[14][1])*(~w6[14][0])) + (window6[15]*(~w6[14][1])*(~w6[14][0]));
           // 01
           channel2[5] = (window6[0]*(~w6[0][1])*(w6[0][0])) + (window6[1]*(~w6[1][1])*(w6[1][0])) + (window6[2]*(~w6[2][1])*(w6[2][0])) + (window6[3]*(~w6[3][1])*(w6[3][0])) + (window6[4]*(~w6[4][1])*(w6[4][0])) + (window6[5]*(~w6[5][1])*(w6[5][0])) + (window6[6]*(~w6[6][1])*(w6[6][0])) + (window6[7]*(~w6[7][1])*(w6[7][0])) + (window6[8]*(~w6[8][1])*(w6[8][0])) + (window6[9]*(~w6[9][1])*(w6[9][0])) + (window6[10]*(~w6[10][1])*(w6[10][0])) + (window6[11]*(~w6[11][1])*(w6[11][0])) +(window6[12]*(~w6[12][1])*(w6[12][0])) + (window6[13]*(~w6[13][1])*(w6[13][0])) + (window6[14]*(~w6[14][1])*(w6[14][0])) + (window6[15]*(~w6[14][1])*(w6[14][0]));
           // 10
           channel3[5] = (window6[0]*(w6[0][1])*(~w6[0][0])) + (window6[1]*(w6[1][1])*(~w6[1][0])) + (window6[2]*(w6[2][1])*(~w6[2][0])) + (window6[3]*(w6[3][1])*(~w6[3][0])) + (window6[4]*(w6[4][1])*(~w6[4][0])) + (window6[5]*(w6[5][1])*(~w6[5][0])) + (window6[6]*(w6[6][1])*(~w6[6][0])) + (window6[7]*(w6[7][1])*(~w6[7][0])) + (window6[8]*(w6[8][1])*(~w6[8][0])) + (window6[9]*(w6[9][1])*(~w6[9][0])) + (window6[10]*(w6[10][1])*(~w6[10][0])) + (window6[11]*(w6[11][1])*(~w6[11][0])) +(window6[12]*(w6[12][1])*(~w6[12][0])) + (window6[13]*(w6[13][1])*(~w6[13][0])) + (window6[14]*(w6[14][1])*(~w6[14][0])) + (window6[15]*(w6[14][1])*(~w6[14][0]));
           // 11
           channel4[5] = (window6[0]*(w6[0][1])*(w6[0][0])) + (window6[1]*(w6[1][1])*(w6[1][0])) + (window6[2]*(w6[2][1])*(w6[2][0])) + (window6[3]*(w6[3][1])*(w6[3][0])) + (window6[4]*(w6[4][1])*(w6[4][0])) + (window6[5]*(w6[5][1])*(w6[5][0])) + (window6[6]*(w6[6][1])*(w6[6][0])) + (window6[7]*(w6[7][1])*(w6[7][0])) + (window6[8]*(w6[8][1])*(w6[8][0])) + (window6[9]*(w6[9][1])*(w6[9][0])) + (window6[10]*(w6[10][1])*(w6[10][0])) + (window6[11]*(w6[11][1])*(w6[11][0])) +(window6[12]*(w6[12][1])*(w6[12][0])) + (window6[13]*(w6[13][1])*(w6[13][0])) + (window6[14]*(w6[14][1])*(w6[14][0])) + (window6[15]*(w6[14][1])*(w6[14][0]));

           // 00
           channel1[6] = (window7[0]*(~w7[0][1])*(~w7[0][0])) + (window7[1]*(~w7[1][1])*(~w7[1][0])) + (window7[2]*(~w7[2][1])*(~w7[2][0])) + (window7[3]*(~w7[3][1])*(~w7[3][0])) + (window7[4]*(~w7[4][1])*(~w7[4][0])) + (window7[5]*(~w7[5][1])*(~w7[5][0])) + (window7[6]*(~w7[6][1])*(~w7[6][0])) + (window7[7]*(~w7[7][1])*(~w7[7][0])) + (window7[8]*(~w7[8][1])*(~w7[8][0])) + (window7[9]*(~w7[9][1])*(~w7[9][0])) + (window7[10]*(~w7[10][1])*(~w7[10][0])) + (window7[11]*(~w7[11][1])*(~w7[11][0])) +(window7[12]*(~w7[12][1])*(~w7[12][0])) + (window7[13]*(~w7[13][1])*(~w7[13][0])) + (window7[14]*(~w7[14][1])*(~w7[14][0])) + (window7[15]*(~w7[14][1])*(~w7[14][0]));
           // 01
           channel2[6] = (window7[0]*(~w7[0][1])*(w7[0][0])) + (window7[1]*(~w7[1][1])*(w7[1][0])) + (window7[2]*(~w7[2][1])*(w7[2][0])) + (window7[3]*(~w7[3][1])*(w7[3][0])) + (window7[4]*(~w7[4][1])*(w7[4][0])) + (window7[5]*(~w7[5][1])*(w7[5][0])) + (window7[6]*(~w7[6][1])*(w7[6][0])) + (window7[7]*(~w7[7][1])*(w7[7][0])) + (window7[8]*(~w7[8][1])*(w7[8][0])) + (window7[9]*(~w7[9][1])*(w7[9][0])) + (window7[10]*(~w7[10][1])*(w7[10][0])) + (window7[11]*(~w7[11][1])*(w7[11][0])) +(window7[12]*(~w7[12][1])*(w7[12][0])) + (window7[13]*(~w7[13][1])*(w7[13][0])) + (window7[14]*(~w7[14][1])*(w7[14][0])) + (window7[15]*(~w7[14][1])*(w7[14][0]));
           // 10
           channel3[6] = (window7[0]*(w7[0][1])*(~w7[0][0])) + (window7[1]*(w7[1][1])*(~w7[1][0])) + (window7[2]*(w7[2][1])*(~w7[2][0])) + (window7[3]*(w7[3][1])*(~w7[3][0])) + (window7[4]*(w7[4][1])*(~w7[4][0])) + (window7[5]*(w7[5][1])*(~w7[5][0])) + (window7[6]*(w7[6][1])*(~w7[6][0])) + (window7[7]*(w7[7][1])*(~w7[7][0])) + (window7[8]*(w7[8][1])*(~w7[8][0])) + (window7[9]*(w7[9][1])*(~w7[9][0])) + (window7[10]*(w7[10][1])*(~w7[10][0])) + (window7[11]*(w7[11][1])*(~w7[11][0])) +(window7[12]*(w7[12][1])*(~w7[12][0])) + (window7[13]*(w7[13][1])*(~w7[13][0])) + (window7[14]*(w7[14][1])*(~w7[14][0])) + (window7[15]*(w7[14][1])*(~w7[14][0]));
           // 11
           channel4[6] = (window7[0]*(w7[0][1])*(w7[0][0])) + (window7[1]*(w7[1][1])*(w7[1][0])) + (window7[2]*(w7[2][1])*(w7[2][0])) + (window7[3]*(w7[3][1])*(w7[3][0])) + (window7[4]*(w7[4][1])*(w7[4][0])) + (window7[5]*(w7[5][1])*(w7[5][0])) + (window7[6]*(w7[6][1])*(w7[6][0])) + (window7[7]*(w7[7][1])*(w7[7][0])) + (window7[8]*(w7[8][1])*(w7[8][0])) + (window7[9]*(w7[9][1])*(w7[9][0])) + (window7[10]*(w7[10][1])*(w7[10][0])) + (window7[11]*(w7[11][1])*(w7[11][0])) +(window7[12]*(w7[12][1])*(w7[12][0])) + (window7[13]*(w7[13][1])*(w7[13][0])) + (window7[14]*(w7[14][1])*(w7[14][0])) + (window7[15]*(w7[14][1])*(w7[14][0]));

           // 00
           channel1[7] = (window8[0]*(~w8[0][1])*(~w8[0][0])) + (window8[1]*(~w8[1][1])*(~w8[1][0])) + (window8[2]*(~w8[2][1])*(~w8[2][0])) + (window8[3]*(~w8[3][1])*(~w8[3][0])) + (window8[4]*(~w8[4][1])*(~w8[4][0])) + (window8[5]*(~w8[5][1])*(~w8[5][0])) + (window8[6]*(~w8[6][1])*(~w8[6][0])) + (window8[7]*(~w8[7][1])*(~w8[7][0])) + (window8[8]*(~w8[8][1])*(~w8[8][0])) + (window8[9]*(~w8[9][1])*(~w8[9][0])) + (window8[10]*(~w8[10][1])*(~w8[10][0])) + (window8[11]*(~w8[11][1])*(~w8[11][0])) +(window8[12]*(~w8[12][1])*(~w8[12][0])) + (window8[13]*(~w8[13][1])*(~w8[13][0])) + (window8[14]*(~w8[14][1])*(~w8[14][0])) + (window8[15]*(~w8[14][1])*(~w8[14][0]));
           // 01
           channel2[7] = (window8[0]*(~w8[0][1])*(w8[0][0])) + (window8[1]*(~w8[1][1])*(w8[1][0])) + (window8[2]*(~w8[2][1])*(w8[2][0])) + (window8[3]*(~w8[3][1])*(w8[3][0])) + (window8[4]*(~w8[4][1])*(w8[4][0])) + (window8[5]*(~w8[5][1])*(w8[5][0])) + (window8[6]*(~w8[6][1])*(w8[6][0])) + (window8[7]*(~w8[7][1])*(w8[7][0])) + (window8[8]*(~w8[8][1])*(w8[8][0])) + (window8[9]*(~w8[9][1])*(w8[9][0])) + (window8[10]*(~w8[10][1])*(w8[10][0])) + (window8[11]*(~w8[11][1])*(w8[11][0])) +(window8[12]*(~w8[12][1])*(w8[12][0])) + (window8[13]*(~w8[13][1])*(w8[13][0])) + (window8[14]*(~w8[14][1])*(w8[14][0])) + (window8[15]*(~w8[14][1])*(w8[14][0]));
           // 10
           channel3[7] = (window8[0]*(w8[0][1])*(~w8[0][0])) + (window8[1]*(w8[1][1])*(~w8[1][0])) + (window8[2]*(w8[2][1])*(~w8[2][0])) + (window8[3]*(w8[3][1])*(~w8[3][0])) + (window8[4]*(w8[4][1])*(~w8[4][0])) + (window8[5]*(w8[5][1])*(~w8[5][0])) + (window8[6]*(w8[6][1])*(~w8[6][0])) + (window8[7]*(w8[7][1])*(~w8[7][0])) + (window8[8]*(w8[8][1])*(~w8[8][0])) + (window8[9]*(w8[9][1])*(~w8[9][0])) + (window8[10]*(w8[10][1])*(~w8[10][0])) + (window8[11]*(w8[11][1])*(~w8[11][0])) +(window8[12]*(w8[12][1])*(~w8[12][0])) + (window8[13]*(w8[13][1])*(~w8[13][0])) + (window8[14]*(w8[14][1])*(~w8[14][0])) + (window8[15]*(w8[14][1])*(~w8[14][0]));
           // 11
           channel4[7] = (window8[0]*(w8[0][1])*(w8[0][0])) + (window8[1]*(w8[1][1])*(w8[1][0])) + (window8[2]*(w8[2][1])*(w8[2][0])) + (window8[3]*(w8[3][1])*(w8[3][0])) + (window8[4]*(w8[4][1])*(w8[4][0])) + (window8[5]*(w8[5][1])*(w8[5][0])) + (window8[6]*(w8[6][1])*(w8[6][0])) + (window8[7]*(w8[7][1])*(w8[7][0])) + (window8[8]*(w8[8][1])*(w8[8][0])) + (window8[9]*(w8[9][1])*(w8[9][0])) + (window8[10]*(w8[10][1])*(w8[10][0])) + (window8[11]*(w8[11][1])*(w8[11][0])) +(window8[12]*(w8[12][1])*(w8[12][0])) + (window8[13]*(w8[13][1])*(w8[13][0])) + (window8[14]*(w8[14][1])*(w8[14][0])) + (window8[15]*(w8[14][1])*(w8[14][0]));

           // 00
           channel1[8] = (window9[0]*(~w9[0][1])*(~w9[0][0])) + (window9[1]*(~w9[1][1])*(~w9[1][0])) + (window9[2]*(~w9[2][1])*(~w9[2][0])) + (window9[3]*(~w9[3][1])*(~w9[3][0])) + (window9[4]*(~w9[4][1])*(~w9[4][0])) + (window9[5]*(~w9[5][1])*(~w9[5][0])) + (window9[6]*(~w9[6][1])*(~w9[6][0])) + (window9[7]*(~w9[7][1])*(~w9[7][0])) + (window9[8]*(~w9[8][1])*(~w9[8][0])) + (window9[9]*(~w9[9][1])*(~w9[9][0])) + (window9[10]*(~w9[10][1])*(~w9[10][0])) + (window9[11]*(~w9[11][1])*(~w9[11][0])) +(window9[12]*(~w9[12][1])*(~w9[12][0])) + (window9[13]*(~w9[13][1])*(~w9[13][0])) + (window9[14]*(~w9[14][1])*(~w9[14][0])) + (window9[15]*(~w9[14][1])*(~w9[14][0]));
           // 01
           channel2[8] = (window9[0]*(~w9[0][1])*(w9[0][0])) + (window9[1]*(~w9[1][1])*(w9[1][0])) + (window9[2]*(~w9[2][1])*(w9[2][0])) + (window9[3]*(~w9[3][1])*(w9[3][0])) + (window9[4]*(~w9[4][1])*(w9[4][0])) + (window9[5]*(~w9[5][1])*(w9[5][0])) + (window9[6]*(~w9[6][1])*(w9[6][0])) + (window9[7]*(~w9[7][1])*(w9[7][0])) + (window9[8]*(~w9[8][1])*(w9[8][0])) + (window9[9]*(~w9[9][1])*(w9[9][0])) + (window9[10]*(~w9[10][1])*(w9[10][0])) + (window9[11]*(~w9[11][1])*(w9[11][0])) +(window9[12]*(~w9[12][1])*(w9[12][0])) + (window9[13]*(~w9[13][1])*(w9[13][0])) + (window9[14]*(~w9[14][1])*(w9[14][0])) + (window9[15]*(~w9[14][1])*(w9[14][0]));
           // 10
           channel3[8] = (window9[0]*(w9[0][1])*(~w9[0][0])) + (window9[1]*(w9[1][1])*(~w9[1][0])) + (window9[2]*(w9[2][1])*(~w9[2][0])) + (window9[3]*(w9[3][1])*(~w9[3][0])) + (window9[4]*(w9[4][1])*(~w9[4][0])) + (window9[5]*(w9[5][1])*(~w9[5][0])) + (window9[6]*(w9[6][1])*(~w9[6][0])) + (window9[7]*(w9[7][1])*(~w9[7][0])) + (window9[8]*(w9[8][1])*(~w9[8][0])) + (window9[9]*(w9[9][1])*(~w9[9][0])) + (window9[10]*(w9[10][1])*(~w9[10][0])) + (window9[11]*(w9[11][1])*(~w9[11][0])) +(window9[12]*(w9[12][1])*(~w9[12][0])) + (window9[13]*(w9[13][1])*(~w9[13][0])) + (window9[14]*(w9[14][1])*(~w9[14][0])) + (window9[15]*(w9[14][1])*(~w9[14][0]));
           // 11
           channel4[8] = (window9[0]*(w9[0][1])*(w9[0][0])) + (window9[1]*(w9[1][1])*(w9[1][0])) + (window9[2]*(w9[2][1])*(w9[2][0])) + (window9[3]*(w9[3][1])*(w9[3][0])) + (window9[4]*(w9[4][1])*(w9[4][0])) + (window9[5]*(w9[5][1])*(w9[5][0])) + (window9[6]*(w9[6][1])*(w9[6][0])) + (window9[7]*(w9[7][1])*(w9[7][0])) + (window9[8]*(w9[8][1])*(w9[8][0])) + (window9[9]*(w9[9][1])*(w9[9][0])) + (window9[10]*(w9[10][1])*(w9[10][0])) + (window9[11]*(w9[11][1])*(w9[11][0])) +(window9[12]*(w9[12][1])*(w9[12][0])) + (window9[13]*(w9[13][1])*(w9[13][0])) + (window9[14]*(w9[14][1])*(w9[14][0])) + (window9[15]*(w9[14][1])*(w9[14][0]));

           // 00
           channel1[9] = (window10[0]*(~w10[0][1])*(~w10[0][0])) + (window10[1]*(~w10[1][1])*(~w10[1][0])) + (window10[2]*(~w10[2][1])*(~w10[2][0])) + (window10[3]*(~w10[3][1])*(~w10[3][0])) + (window10[4]*(~w10[4][1])*(~w10[4][0])) + (window10[5]*(~w10[5][1])*(~w10[5][0])) + (window10[6]*(~w10[6][1])*(~w10[6][0])) + (window10[7]*(~w10[7][1])*(~w10[7][0])) + (window10[8]*(~w10[8][1])*(~w10[8][0])) + (window10[9]*(~w10[9][1])*(~w10[9][0])) + (window10[10]*(~w10[10][1])*(~w10[10][0])) + (window10[11]*(~w10[11][1])*(~w10[11][0])) +(window10[12]*(~w10[12][1])*(~w10[12][0])) + (window10[13]*(~w10[13][1])*(~w10[13][0])) + (window10[14]*(~w10[14][1])*(~w10[14][0])) + (window10[15]*(~w10[14][1])*(~w10[14][0]));
           // 01
           channel2[9] = (window10[0]*(~w10[0][1])*(w10[0][0])) + (window10[1]*(~w10[1][1])*(w10[1][0])) + (window10[2]*(~w10[2][1])*(w10[2][0])) + (window10[3]*(~w10[3][1])*(w10[3][0])) + (window10[4]*(~w10[4][1])*(w10[4][0])) + (window10[5]*(~w10[5][1])*(w10[5][0])) + (window10[6]*(~w10[6][1])*(w10[6][0])) + (window10[7]*(~w10[7][1])*(w10[7][0])) + (window10[8]*(~w10[8][1])*(w10[8][0])) + (window10[9]*(~w10[9][1])*(w10[9][0])) + (window10[10]*(~w10[10][1])*(w10[10][0])) + (window10[11]*(~w10[11][1])*(w10[11][0])) +(window10[12]*(~w10[12][1])*(w10[12][0])) + (window10[13]*(~w10[13][1])*(w10[13][0])) + (window10[14]*(~w10[14][1])*(w10[14][0])) + (window10[15]*(~w10[14][1])*(w10[14][0]));
           // 10
           channel3[9] = (window10[0]*(w10[0][1])*(~w10[0][0])) + (window10[1]*(w10[1][1])*(~w10[1][0])) + (window10[2]*(w10[2][1])*(~w10[2][0])) + (window10[3]*(w10[3][1])*(~w10[3][0])) + (window10[4]*(w10[4][1])*(~w10[4][0])) + (window10[5]*(w10[5][1])*(~w10[5][0])) + (window10[6]*(w10[6][1])*(~w10[6][0])) + (window10[7]*(w10[7][1])*(~w10[7][0])) + (window10[8]*(w10[8][1])*(~w10[8][0])) + (window10[9]*(w10[9][1])*(~w10[9][0])) + (window10[10]*(w10[10][1])*(~w10[10][0])) + (window10[11]*(w10[11][1])*(~w10[11][0])) +(window10[12]*(w10[12][1])*(~w10[12][0])) + (window10[13]*(w10[13][1])*(~w10[13][0])) + (window10[14]*(w10[14][1])*(~w10[14][0])) + (window10[15]*(w10[14][1])*(~w10[14][0]));
           // 11
           channel4[9] = (window10[0]*(w10[0][1])*(w10[0][0])) + (window10[1]*(w10[1][1])*(w10[1][0])) + (window10[2]*(w10[2][1])*(w10[2][0])) + (window10[3]*(w10[3][1])*(w10[3][0])) + (window10[4]*(w10[4][1])*(w10[4][0])) + (window10[5]*(w10[5][1])*(w10[5][0])) + (window10[6]*(w10[6][1])*(w10[6][0])) + (window10[7]*(w10[7][1])*(w10[7][0])) + (window10[8]*(w10[8][1])*(w10[8][0])) + (window10[9]*(w10[9][1])*(w10[9][0])) + (window10[10]*(w10[10][1])*(w10[10][0])) + (window10[11]*(w10[11][1])*(w10[11][0])) +(window10[12]*(w10[12][1])*(w10[12][0])) + (window10[13]*(w10[13][1])*(w10[13][0])) + (window10[14]*(w10[14][1])*(w10[14][0])) + (window10[15]*(w10[14][1])*(w10[14][0]));

           // 00
           channel1[10] = (window11[0]*(~w11[0][1])*(~w11[0][0])) + (window11[1]*(~w11[1][1])*(~w11[1][0])) + (window11[2]*(~w11[2][1])*(~w11[2][0])) + (window11[3]*(~w11[3][1])*(~w11[3][0])) + (window11[4]*(~w11[4][1])*(~w11[4][0])) + (window11[5]*(~w11[5][1])*(~w11[5][0])) + (window11[6]*(~w11[6][1])*(~w11[6][0])) + (window11[7]*(~w11[7][1])*(~w11[7][0])) + (window11[8]*(~w11[8][1])*(~w11[8][0])) + (window11[9]*(~w11[9][1])*(~w11[9][0])) + (window11[10]*(~w11[10][1])*(~w11[10][0])) + (window11[11]*(~w11[11][1])*(~w11[11][0])) +(window11[12]*(~w11[12][1])*(~w11[12][0])) + (window11[13]*(~w11[13][1])*(~w11[13][0])) + (window11[14]*(~w11[14][1])*(~w11[14][0])) + (window11[15]*(~w11[14][1])*(~w11[14][0]));
           // 01
           channel2[10] = (window11[0]*(~w11[0][1])*(w11[0][0])) + (window11[1]*(~w11[1][1])*(w11[1][0])) + (window11[2]*(~w11[2][1])*(w11[2][0])) + (window11[3]*(~w11[3][1])*(w11[3][0])) + (window11[4]*(~w11[4][1])*(w11[4][0])) + (window11[5]*(~w11[5][1])*(w11[5][0])) + (window11[6]*(~w11[6][1])*(w11[6][0])) + (window11[7]*(~w11[7][1])*(w11[7][0])) + (window11[8]*(~w11[8][1])*(w11[8][0])) + (window11[9]*(~w11[9][1])*(w11[9][0])) + (window11[10]*(~w11[10][1])*(w11[10][0])) + (window11[11]*(~w11[11][1])*(w11[11][0])) +(window11[12]*(~w11[12][1])*(w11[12][0])) + (window11[13]*(~w11[13][1])*(w11[13][0])) + (window11[14]*(~w11[14][1])*(w11[14][0])) + (window11[15]*(~w11[14][1])*(w11[14][0]));
           // 10
           channel3[10] = (window11[0]*(w11[0][1])*(~w11[0][0])) + (window11[1]*(w11[1][1])*(~w11[1][0])) + (window11[2]*(w11[2][1])*(~w11[2][0])) + (window11[3]*(w11[3][1])*(~w11[3][0])) + (window11[4]*(w11[4][1])*(~w11[4][0])) + (window11[5]*(w11[5][1])*(~w11[5][0])) + (window11[6]*(w11[6][1])*(~w11[6][0])) + (window11[7]*(w11[7][1])*(~w11[7][0])) + (window11[8]*(w11[8][1])*(~w11[8][0])) + (window11[9]*(w11[9][1])*(~w11[9][0])) + (window11[10]*(w11[10][1])*(~w11[10][0])) + (window11[11]*(w11[11][1])*(~w11[11][0])) +(window11[12]*(w11[12][1])*(~w11[12][0])) + (window11[13]*(w11[13][1])*(~w11[13][0])) + (window11[14]*(w11[14][1])*(~w11[14][0])) + (window11[15]*(w11[14][1])*(~w11[14][0]));
           // 11
           channel4[10] = (window11[0]*(w11[0][1])*(w11[0][0])) + (window11[1]*(w11[1][1])*(w11[1][0])) + (window11[2]*(w11[2][1])*(w11[2][0])) + (window11[3]*(w11[3][1])*(w11[3][0])) + (window11[4]*(w11[4][1])*(w11[4][0])) + (window11[5]*(w11[5][1])*(w11[5][0])) + (window11[6]*(w11[6][1])*(w11[6][0])) + (window11[7]*(w11[7][1])*(w11[7][0])) + (window11[8]*(w11[8][1])*(w11[8][0])) + (window11[9]*(w11[9][1])*(w11[9][0])) + (window11[10]*(w11[10][1])*(w11[10][0])) + (window11[11]*(w11[11][1])*(w11[11][0])) +(window11[12]*(w11[12][1])*(w11[12][0])) + (window11[13]*(w11[13][1])*(w11[13][0])) + (window11[14]*(w11[14][1])*(w11[14][0])) + (window11[15]*(w11[14][1])*(w11[14][0]));

           // 00
           channel1[11] = (window12[0]*(~w12[0][1])*(~w12[0][0])) + (window12[1]*(~w12[1][1])*(~w12[1][0])) + (window12[2]*(~w12[2][1])*(~w12[2][0])) + (window12[3]*(~w12[3][1])*(~w12[3][0])) + (window12[4]*(~w12[4][1])*(~w12[4][0])) + (window12[5]*(~w12[5][1])*(~w12[5][0])) + (window12[6]*(~w12[6][1])*(~w12[6][0])) + (window12[7]*(~w12[7][1])*(~w12[7][0])) + (window12[8]*(~w12[8][1])*(~w12[8][0])) + (window12[9]*(~w12[9][1])*(~w12[9][0])) + (window12[10]*(~w12[10][1])*(~w12[10][0])) + (window12[11]*(~w12[11][1])*(~w12[11][0])) +(window12[12]*(~w12[12][1])*(~w12[12][0])) + (window12[13]*(~w12[13][1])*(~w12[13][0])) + (window12[14]*(~w12[14][1])*(~w12[14][0])) + (window12[15]*(~w12[14][1])*(~w12[14][0]));
           // 01
           channel2[11] = (window12[0]*(~w12[0][1])*(w12[0][0])) + (window12[1]*(~w12[1][1])*(w12[1][0])) + (window12[2]*(~w12[2][1])*(w12[2][0])) + (window12[3]*(~w12[3][1])*(w12[3][0])) + (window12[4]*(~w12[4][1])*(w12[4][0])) + (window12[5]*(~w12[5][1])*(w12[5][0])) + (window12[6]*(~w12[6][1])*(w12[6][0])) + (window12[7]*(~w12[7][1])*(w12[7][0])) + (window12[8]*(~w12[8][1])*(w12[8][0])) + (window12[9]*(~w12[9][1])*(w12[9][0])) + (window12[10]*(~w12[10][1])*(w12[10][0])) + (window12[11]*(~w12[11][1])*(w12[11][0])) +(window12[12]*(~w12[12][1])*(w12[12][0])) + (window12[13]*(~w12[13][1])*(w12[13][0])) + (window12[14]*(~w12[14][1])*(w12[14][0])) + (window12[15]*(~w12[14][1])*(w12[14][0]));
           // 10
           channel3[11] = (window12[0]*(w12[0][1])*(~w12[0][0])) + (window12[1]*(w12[1][1])*(~w12[1][0])) + (window12[2]*(w12[2][1])*(~w12[2][0])) + (window12[3]*(w12[3][1])*(~w12[3][0])) + (window12[4]*(w12[4][1])*(~w12[4][0])) + (window12[5]*(w12[5][1])*(~w12[5][0])) + (window12[6]*(w12[6][1])*(~w12[6][0])) + (window12[7]*(w12[7][1])*(~w12[7][0])) + (window12[8]*(w12[8][1])*(~w12[8][0])) + (window12[9]*(w12[9][1])*(~w12[9][0])) + (window12[10]*(w12[10][1])*(~w12[10][0])) + (window12[11]*(w12[11][1])*(~w12[11][0])) +(window12[12]*(w12[12][1])*(~w12[12][0])) + (window12[13]*(w12[13][1])*(~w12[13][0])) + (window12[14]*(w12[14][1])*(~w12[14][0])) + (window12[15]*(w12[14][1])*(~w12[14][0]));
           // 11
           channel4[11] = (window12[0]*(w12[0][1])*(w12[0][0])) + (window12[1]*(w12[1][1])*(w12[1][0])) + (window12[2]*(w12[2][1])*(w12[2][0])) + (window12[3]*(w12[3][1])*(w12[3][0])) + (window12[4]*(w12[4][1])*(w12[4][0])) + (window12[5]*(w12[5][1])*(w12[5][0])) + (window12[6]*(w12[6][1])*(w12[6][0])) + (window12[7]*(w12[7][1])*(w12[7][0])) + (window12[8]*(w12[8][1])*(w12[8][0])) + (window12[9]*(w12[9][1])*(w12[9][0])) + (window12[10]*(w12[10][1])*(w12[10][0])) + (window12[11]*(w12[11][1])*(w12[11][0])) +(window12[12]*(w12[12][1])*(w12[12][0])) + (window12[13]*(w12[13][1])*(w12[13][0])) + (window12[14]*(w12[14][1])*(w12[14][0])) + (window12[15]*(w12[14][1])*(w12[14][0]));

           // 00
           channel1[12] = (window13[0]*(~w13[0][1])*(~w13[0][0])) + (window13[1]*(~w13[1][1])*(~w13[1][0])) + (window13[2]*(~w13[2][1])*(~w13[2][0])) + (window13[3]*(~w13[3][1])*(~w13[3][0])) + (window13[4]*(~w13[4][1])*(~w13[4][0])) + (window13[5]*(~w13[5][1])*(~w13[5][0])) + (window13[6]*(~w13[6][1])*(~w13[6][0])) + (window13[7]*(~w13[7][1])*(~w13[7][0])) + (window13[8]*(~w13[8][1])*(~w13[8][0])) + (window13[9]*(~w13[9][1])*(~w13[9][0])) + (window13[10]*(~w13[10][1])*(~w13[10][0])) + (window13[11]*(~w13[11][1])*(~w13[11][0])) +(window13[12]*(~w13[12][1])*(~w13[12][0])) + (window13[13]*(~w13[13][1])*(~w13[13][0])) + (window13[14]*(~w13[14][1])*(~w13[14][0])) + (window13[15]*(~w13[14][1])*(~w13[14][0]));
           // 01
           channel2[12] = (window13[0]*(~w13[0][1])*(w13[0][0])) + (window13[1]*(~w13[1][1])*(w13[1][0])) + (window13[2]*(~w13[2][1])*(w13[2][0])) + (window13[3]*(~w13[3][1])*(w13[3][0])) + (window13[4]*(~w13[4][1])*(w13[4][0])) + (window13[5]*(~w13[5][1])*(w13[5][0])) + (window13[6]*(~w13[6][1])*(w13[6][0])) + (window13[7]*(~w13[7][1])*(w13[7][0])) + (window13[8]*(~w13[8][1])*(w13[8][0])) + (window13[9]*(~w13[9][1])*(w13[9][0])) + (window13[10]*(~w13[10][1])*(w13[10][0])) + (window13[11]*(~w13[11][1])*(w13[11][0])) +(window13[12]*(~w13[12][1])*(w13[12][0])) + (window13[13]*(~w13[13][1])*(w13[13][0])) + (window13[14]*(~w13[14][1])*(w13[14][0])) + (window13[15]*(~w13[14][1])*(w13[14][0]));
           // 10
           channel3[12] = (window13[0]*(w13[0][1])*(~w13[0][0])) + (window13[1]*(w13[1][1])*(~w13[1][0])) + (window13[2]*(w13[2][1])*(~w13[2][0])) + (window13[3]*(w13[3][1])*(~w13[3][0])) + (window13[4]*(w13[4][1])*(~w13[4][0])) + (window13[5]*(w13[5][1])*(~w13[5][0])) + (window13[6]*(w13[6][1])*(~w13[6][0])) + (window13[7]*(w13[7][1])*(~w13[7][0])) + (window13[8]*(w13[8][1])*(~w13[8][0])) + (window13[9]*(w13[9][1])*(~w13[9][0])) + (window13[10]*(w13[10][1])*(~w13[10][0])) + (window13[11]*(w13[11][1])*(~w13[11][0])) +(window13[12]*(w13[12][1])*(~w13[12][0])) + (window13[13]*(w13[13][1])*(~w13[13][0])) + (window13[14]*(w13[14][1])*(~w13[14][0])) + (window13[15]*(w13[14][1])*(~w13[14][0]));
           // 11
           channel4[12] = (window13[0]*(w13[0][1])*(w13[0][0])) + (window13[1]*(w13[1][1])*(w13[1][0])) + (window13[2]*(w13[2][1])*(w13[2][0])) + (window13[3]*(w13[3][1])*(w13[3][0])) + (window13[4]*(w13[4][1])*(w13[4][0])) + (window13[5]*(w13[5][1])*(w13[5][0])) + (window13[6]*(w13[6][1])*(w13[6][0])) + (window13[7]*(w13[7][1])*(w13[7][0])) + (window13[8]*(w13[8][1])*(w13[8][0])) + (window13[9]*(w13[9][1])*(w13[9][0])) + (window13[10]*(w13[10][1])*(w13[10][0])) + (window13[11]*(w13[11][1])*(w13[11][0])) +(window13[12]*(w13[12][1])*(w13[12][0])) + (window13[13]*(w13[13][1])*(w13[13][0])) + (window13[14]*(w13[14][1])*(w13[14][0])) + (window13[15]*(w13[14][1])*(w13[14][0]));

           // 00
           channel1[13] = (window14[0]*(~w14[0][1])*(~w14[0][0])) + (window14[1]*(~w14[1][1])*(~w14[1][0])) + (window14[2]*(~w14[2][1])*(~w14[2][0])) + (window14[3]*(~w14[3][1])*(~w14[3][0])) + (window14[4]*(~w14[4][1])*(~w14[4][0])) + (window14[5]*(~w14[5][1])*(~w14[5][0])) + (window14[6]*(~w14[6][1])*(~w14[6][0])) + (window14[7]*(~w14[7][1])*(~w14[7][0])) + (window14[8]*(~w14[8][1])*(~w14[8][0])) + (window14[9]*(~w14[9][1])*(~w14[9][0])) + (window14[10]*(~w14[10][1])*(~w14[10][0])) + (window14[11]*(~w14[11][1])*(~w14[11][0])) +(window14[12]*(~w14[12][1])*(~w14[12][0])) + (window14[13]*(~w14[13][1])*(~w14[13][0])) + (window14[14]*(~w14[14][1])*(~w14[14][0])) + (window14[15]*(~w14[14][1])*(~w14[14][0]));
           // 01
           channel2[13] = (window14[0]*(~w14[0][1])*(w14[0][0])) + (window14[1]*(~w14[1][1])*(w14[1][0])) + (window14[2]*(~w14[2][1])*(w14[2][0])) + (window14[3]*(~w14[3][1])*(w14[3][0])) + (window14[4]*(~w14[4][1])*(w14[4][0])) + (window14[5]*(~w14[5][1])*(w14[5][0])) + (window14[6]*(~w14[6][1])*(w14[6][0])) + (window14[7]*(~w14[7][1])*(w14[7][0])) + (window14[8]*(~w14[8][1])*(w14[8][0])) + (window14[9]*(~w14[9][1])*(w14[9][0])) + (window14[10]*(~w14[10][1])*(w14[10][0])) + (window14[11]*(~w14[11][1])*(w14[11][0])) +(window14[12]*(~w14[12][1])*(w14[12][0])) + (window14[13]*(~w14[13][1])*(w14[13][0])) + (window14[14]*(~w14[14][1])*(w14[14][0])) + (window14[15]*(~w14[14][1])*(w14[14][0]));
           // 10
           channel3[13] = (window14[0]*(w14[0][1])*(~w14[0][0])) + (window14[1]*(w14[1][1])*(~w14[1][0])) + (window14[2]*(w14[2][1])*(~w14[2][0])) + (window14[3]*(w14[3][1])*(~w14[3][0])) + (window14[4]*(w14[4][1])*(~w14[4][0])) + (window14[5]*(w14[5][1])*(~w14[5][0])) + (window14[6]*(w14[6][1])*(~w14[6][0])) + (window14[7]*(w14[7][1])*(~w14[7][0])) + (window14[8]*(w14[8][1])*(~w14[8][0])) + (window14[9]*(w14[9][1])*(~w14[9][0])) + (window14[10]*(w14[10][1])*(~w14[10][0])) + (window14[11]*(w14[11][1])*(~w14[11][0])) +(window14[12]*(w14[12][1])*(~w14[12][0])) + (window14[13]*(w14[13][1])*(~w14[13][0])) + (window14[14]*(w14[14][1])*(~w14[14][0])) + (window14[15]*(w14[14][1])*(~w14[14][0]));
           // 11
           channel4[13] = (window14[0]*(w14[0][1])*(w14[0][0])) + (window14[1]*(w14[1][1])*(w14[1][0])) + (window14[2]*(w14[2][1])*(w14[2][0])) + (window14[3]*(w14[3][1])*(w14[3][0])) + (window14[4]*(w14[4][1])*(w14[4][0])) + (window14[5]*(w14[5][1])*(w14[5][0])) + (window14[6]*(w14[6][1])*(w14[6][0])) + (window14[7]*(w14[7][1])*(w14[7][0])) + (window14[8]*(w14[8][1])*(w14[8][0])) + (window14[9]*(w14[9][1])*(w14[9][0])) + (window14[10]*(w14[10][1])*(w14[10][0])) + (window14[11]*(w14[11][1])*(w14[11][0])) +(window14[12]*(w14[12][1])*(w14[12][0])) + (window14[13]*(w14[13][1])*(w14[13][0])) + (window14[14]*(w14[14][1])*(w14[14][0])) + (window14[15]*(w14[14][1])*(w14[14][0]));

           // 00
           channel1[14] = (window15[0]*(~w15[0][1])*(~w15[0][0])) + (window15[1]*(~w15[1][1])*(~w15[1][0])) + (window15[2]*(~w15[2][1])*(~w15[2][0])) + (window15[3]*(~w15[3][1])*(~w15[3][0])) + (window15[4]*(~w15[4][1])*(~w15[4][0])) + (window15[5]*(~w15[5][1])*(~w15[5][0])) + (window15[6]*(~w15[6][1])*(~w15[6][0])) + (window15[7]*(~w15[7][1])*(~w15[7][0])) + (window15[8]*(~w15[8][1])*(~w15[8][0])) + (window15[9]*(~w15[9][1])*(~w15[9][0])) + (window15[10]*(~w15[10][1])*(~w15[10][0])) + (window15[11]*(~w15[11][1])*(~w15[11][0])) +(window15[12]*(~w15[12][1])*(~w15[12][0])) + (window15[13]*(~w15[13][1])*(~w15[13][0])) + (window15[14]*(~w15[14][1])*(~w15[14][0])) + (window15[15]*(~w15[14][1])*(~w15[14][0]));
           // 01
           channel2[14] = (window15[0]*(~w15[0][1])*(w15[0][0])) + (window15[1]*(~w15[1][1])*(w15[1][0])) + (window15[2]*(~w15[2][1])*(w15[2][0])) + (window15[3]*(~w15[3][1])*(w15[3][0])) + (window15[4]*(~w15[4][1])*(w15[4][0])) + (window15[5]*(~w15[5][1])*(w15[5][0])) + (window15[6]*(~w15[6][1])*(w15[6][0])) + (window15[7]*(~w15[7][1])*(w15[7][0])) + (window15[8]*(~w15[8][1])*(w15[8][0])) + (window15[9]*(~w15[9][1])*(w15[9][0])) + (window15[10]*(~w15[10][1])*(w15[10][0])) + (window15[11]*(~w15[11][1])*(w15[11][0])) +(window15[12]*(~w15[12][1])*(w15[12][0])) + (window15[13]*(~w15[13][1])*(w15[13][0])) + (window15[14]*(~w15[14][1])*(w15[14][0])) + (window15[15]*(~w15[14][1])*(w15[14][0]));
           // 10
           channel3[14] = (window15[0]*(w15[0][1])*(~w15[0][0])) + (window15[1]*(w15[1][1])*(~w15[1][0])) + (window15[2]*(w15[2][1])*(~w15[2][0])) + (window15[3]*(w15[3][1])*(~w15[3][0])) + (window15[4]*(w15[4][1])*(~w15[4][0])) + (window15[5]*(w15[5][1])*(~w15[5][0])) + (window15[6]*(w15[6][1])*(~w15[6][0])) + (window15[7]*(w15[7][1])*(~w15[7][0])) + (window15[8]*(w15[8][1])*(~w15[8][0])) + (window15[9]*(w15[9][1])*(~w15[9][0])) + (window15[10]*(w15[10][1])*(~w15[10][0])) + (window15[11]*(w15[11][1])*(~w15[11][0])) +(window15[12]*(w15[12][1])*(~w15[12][0])) + (window15[13]*(w15[13][1])*(~w15[13][0])) + (window15[14]*(w15[14][1])*(~w15[14][0])) + (window15[15]*(w15[14][1])*(~w15[14][0]));
           // 11
           channel4[14] = (window15[0]*(w15[0][1])*(w15[0][0])) + (window15[1]*(w15[1][1])*(w15[1][0])) + (window15[2]*(w15[2][1])*(w15[2][0])) + (window15[3]*(w15[3][1])*(w15[3][0])) + (window15[4]*(w15[4][1])*(w15[4][0])) + (window15[5]*(w15[5][1])*(w15[5][0])) + (window15[6]*(w15[6][1])*(w15[6][0])) + (window15[7]*(w15[7][1])*(w15[7][0])) + (window15[8]*(w15[8][1])*(w15[8][0])) + (window15[9]*(w15[9][1])*(w15[9][0])) + (window15[10]*(w15[10][1])*(w15[10][0])) + (window15[11]*(w15[11][1])*(w15[11][0])) +(window15[12]*(w15[12][1])*(w15[12][0])) + (window15[13]*(w15[13][1])*(w15[13][0])) + (window15[14]*(w15[14][1])*(w15[14][0])) + (window15[15]*(w15[14][1])*(w15[14][0]));

           // 00
           channel1[15] = (window16[0]*(~w16[0][1])*(~w16[0][0])) + (window16[1]*(~w16[1][1])*(~w16[1][0])) + (window16[2]*(~w16[2][1])*(~w16[2][0])) + (window16[3]*(~w16[3][1])*(~w16[3][0])) + (window16[4]*(~w16[4][1])*(~w16[4][0])) + (window16[5]*(~w16[5][1])*(~w16[5][0])) + (window16[6]*(~w16[6][1])*(~w16[6][0])) + (window16[7]*(~w16[7][1])*(~w16[7][0])) + (window16[8]*(~w16[8][1])*(~w16[8][0])) + (window16[9]*(~w16[9][1])*(~w16[9][0])) + (window16[10]*(~w16[10][1])*(~w16[10][0])) + (window16[11]*(~w16[11][1])*(~w16[11][0])) +(window16[12]*(~w16[12][1])*(~w16[12][0])) + (window16[13]*(~w16[13][1])*(~w16[13][0])) + (window16[14]*(~w16[14][1])*(~w16[14][0])) + (window16[15]*(~w16[14][1])*(~w16[14][0]));
           // 01
           channel2[15] = (window16[0]*(~w16[0][1])*(w16[0][0])) + (window16[1]*(~w16[1][1])*(w16[1][0])) + (window16[2]*(~w16[2][1])*(w16[2][0])) + (window16[3]*(~w16[3][1])*(w16[3][0])) + (window16[4]*(~w16[4][1])*(w16[4][0])) + (window16[5]*(~w16[5][1])*(w16[5][0])) + (window16[6]*(~w16[6][1])*(w16[6][0])) + (window16[7]*(~w16[7][1])*(w16[7][0])) + (window16[8]*(~w16[8][1])*(w16[8][0])) + (window16[9]*(~w16[9][1])*(w16[9][0])) + (window16[10]*(~w16[10][1])*(w16[10][0])) + (window16[11]*(~w16[11][1])*(w16[11][0])) +(window16[12]*(~w16[12][1])*(w16[12][0])) + (window16[13]*(~w16[13][1])*(w16[13][0])) + (window16[14]*(~w16[14][1])*(w16[14][0])) + (window16[15]*(~w16[14][1])*(w16[14][0]));
           // 10
           channel3[15] = (window16[0]*(w16[0][1])*(~w16[0][0])) + (window16[1]*(w16[1][1])*(~w16[1][0])) + (window16[2]*(w16[2][1])*(~w16[2][0])) + (window16[3]*(w16[3][1])*(~w16[3][0])) + (window16[4]*(w16[4][1])*(~w16[4][0])) + (window16[5]*(w16[5][1])*(~w16[5][0])) + (window16[6]*(w16[6][1])*(~w16[6][0])) + (window16[7]*(w16[7][1])*(~w16[7][0])) + (window16[8]*(w16[8][1])*(~w16[8][0])) + (window16[9]*(w16[9][1])*(~w16[9][0])) + (window16[10]*(w16[10][1])*(~w16[10][0])) + (window16[11]*(w16[11][1])*(~w16[11][0])) +(window16[12]*(w16[12][1])*(~w16[12][0])) + (window16[13]*(w16[13][1])*(~w16[13][0])) + (window16[14]*(w16[14][1])*(~w16[14][0])) + (window16[15]*(w16[14][1])*(~w16[14][0]));
           // 11
           channel4[15] = (window16[0]*(w16[0][1])*(w16[0][0])) + (window16[1]*(w16[1][1])*(w16[1][0])) + (window16[2]*(w16[2][1])*(w16[2][0])) + (window16[3]*(w16[3][1])*(w16[3][0])) + (window16[4]*(w16[4][1])*(w16[4][0])) + (window16[5]*(w16[5][1])*(w16[5][0])) + (window16[6]*(w16[6][1])*(w16[6][0])) + (window16[7]*(w16[7][1])*(w16[7][0])) + (window16[8]*(w16[8][1])*(w16[8][0])) + (window16[9]*(w16[9][1])*(w16[9][0])) + (window16[10]*(w16[10][1])*(w16[10][0])) + (window16[11]*(w16[11][1])*(w16[11][0])) +(window16[12]*(w16[12][1])*(w16[12][0])) + (window16[13]*(w16[13][1])*(w16[13][0])) + (window16[14]*(w16[14][1])*(w16[14][0])) + (window16[15]*(w16[14][1])*(w16[14][0]));

           NS = COMPUTE;
          end
 COMPUTE: begin
           descriptor_1 = channel1[0] + channel1[1] + channel1[2] + channel1[3] + channel1[4] + channel1[5] + channel1[6] + channel1[7] + channel1[8] + channel1[9] + channel1[10] + channel1[11] + channel1[12] + channel1[13] + channel1[14] + channel1[15];
           descriptor_2 = channel2[0] + channel2[1] + channel2[2] + channel2[3] + channel2[4] + channel2[5] + channel2[6] + channel2[7] + channel2[8] + channel2[9] + channel2[10] + channel2[11] + channel2[12] + channel2[13] + channel2[14] + channel2[15];
           descriptor_3 = channel3[0] + channel3[1] + channel3[2] + channel3[3] + channel3[4] + channel3[5] + channel3[6] + channel3[7] + channel3[8] + channel3[9] + channel3[10] + channel3[11] + channel3[12] + channel3[13] + channel3[14] + channel3[15];
           descriptor_4 = channel4[0] + channel4[1] + channel4[2] + channel4[3] + channel4[4] + channel4[5] + channel4[6] + channel4[7] + channel4[8] + channel4[9] + channel4[10] + channel4[11] + channel4[12] + channel4[13] + channel4[14] + channel4[15];

           NS = ASSIGN;
          end
 endcase
end
assign output_valid = (PS == COMPUTE) ? 1'b1 : 1'b0;
assign keypoint = (PS == COMPUTE) ? k : 32'hzzzzzzzz;
assign descriptor_channel_1 = (PS == COMPUTE) ? descriptor_1 : 16'hzzzz;
assign descriptor_channel_2 = (PS == COMPUTE) ? descriptor_2 : 16'hzzzz;
assign descriptor_channel_3 = (PS == COMPUTE) ? descriptor_3 : 16'hzzzz;
assign descriptor_channel_4 = (PS == COMPUTE) ? descriptor_4 : 16'hzzzz;
assign done = (count == limit-1) ? 1'b1 : 1'b0;
endmodule
